* Extracted by KLayout with SG13G2 LVS runset on : 12/02/2026 15:34

.SUBCKT T_gate gnd vdd Control Vout Vin \!Control
M$1 Vin Control Vout gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$2 Vin \!Control Vout vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
.ENDS T_gate
