** sch_path: /home/designer/shared/IHP-AnalogAcademy/modules/module_3_8_bit_SAR_ADC/part_5_analog_layout/switch_array/schematic/T_gate_switch.sch
.subckt T_gate_switch Vo Control vdd vref gnd
*.PININFO Vo:B Control:B vdd:B vref:B gnd:B
x12 net1 gnd Vo gnd Control vdd T_gate
x14 Control vref Vo gnd net1 vdd T_gate
x13 vdd Control net1 gnd inverter
.ends

* expanding   symbol:  T_gate.sym # of pins=6
** sym_path: /home/designer/shared/IHP-AnalogAcademy/modules/module_3_8_bit_SAR_ADC/part_5_analog_layout/switch_array/schematic/T_gate.sym
** sch_path: /home/designer/shared/IHP-AnalogAcademy/modules/module_3_8_bit_SAR_ADC/part_5_analog_layout/switch_array/schematic/T_gate.sch
.subckt T_gate !Control Vin Vout gnd Control vdd
*.PININFO Vout:B Vin:B !Control:B Control:B gnd:B vdd:B
M1 Vin Control Vout gnd sg13_lv_nmos w=1u l=0.13u ng=1 m=1
M2 Vin !Control Vout vdd sg13_lv_pmos w=2u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/designer/shared/IHP-AnalogAcademy/modules/module_3_8_bit_SAR_ADC/part_5_analog_layout/switch_array/schematic/inverter.sym
** sch_path: /home/designer/shared/IHP-AnalogAcademy/modules/module_3_8_bit_SAR_ADC/part_5_analog_layout/switch_array/schematic/inverter.sch
.subckt inverter vdd vi vo gnd
*.PININFO vi:B vo:B gnd:B vdd:B
M5 vo vi vdd vdd sg13_lv_pmos w=800n l=130n ng=1 m=1
M7 vo vi gnd gnd sg13_lv_nmos w=400n l=130n ng=1 m=1
.ends

