** sch_path: /home/designer/shared/IHP-AnalogAcademy/modules/module_3_8_bit_SAR_ADC/part_5_analog_layout/switch_array/schematic/inverter.sch
.subckt inverter vdd vi vo gnd
*.PININFO vi:B vo:B gnd:B vdd:B
M5 vo vi vdd vdd sg13_lv_pmos w=800n l=130n ng=1 m=1
M7 vo vi gnd gnd sg13_lv_nmos w=400n l=130n ng=1 m=1
.ends
