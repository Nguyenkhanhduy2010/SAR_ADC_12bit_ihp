* Extracted by KLayout with SG13G2 LVS runset on : 26/02/2026 12:18

.SUBCKT CDAC C_MSB vo C6 C5 vref C4 C1 C3 C2
C$1 \$3 \$2 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=40
C$14 vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=64
C$41 vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=32
C$56 vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=16
C$60 vo vref cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$69 vo C4 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=8
C$72 vo C1 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$82 vo C3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=4
C$83 vo C2 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=2
.ENDS CDAC
