* Extracted by KLayout with SG13G2 LVS runset on : 26/02/2026 08:15

.SUBCKT DIFF_COMPARATOR clk gnd vdd vbias out\x2d out+ V+ V\x2d
M$1 gnd gnd gnd \$1 sg13_lv_nmos L=0.2u W=16u AS=4.24p AD=4.24p PS=26.12u
+ PD=26.12u
M$2 gnd clk \$8 \$1 sg13_lv_nmos L=0.2u W=4u AS=0.76p AD=1.44p PS=4.38u PD=4.72u
M$3 \$8 \$9 gnd \$1 sg13_lv_nmos L=0.2u W=4u AS=1.44p AD=0.76p PS=4.72u PD=4.38u
M$6 gnd \$8 \$9 \$1 sg13_lv_nmos L=0.2u W=4u AS=0.76p AD=1.44p PS=4.38u PD=4.72u
M$7 \$9 clk gnd \$1 sg13_lv_nmos L=0.2u W=4u AS=1.44p AD=0.76p PS=4.72u PD=4.38u
M$9 out\x2d \$8 gnd \$1 sg13_lv_nmos L=0.2u W=4u AS=1.06p AD=1.06p PS=7.06u
+ PD=7.06u
M$11 out+ \$9 gnd \$1 sg13_lv_nmos L=0.2u W=4u AS=1.06p AD=1.06p PS=7.06u
+ PD=7.06u
M$13 \$7 vbias vdd \$5 sg13_lv_pmos L=0.3u W=18u AS=4.095p AD=4.095p PS=24.32u
+ PD=24.32u
M$17 \$26 clk \$7 \$5 sg13_lv_pmos L=0.3u W=18u AS=4.095p AD=4.095p PS=24.32u
+ PD=24.32u
M$21 out\x2d \$8 vdd \$5 sg13_lv_pmos L=0.2u W=8u AS=2.12p AD=2.12p PS=13.06u
+ PD=13.06u
M$23 out+ \$9 vdd \$5 sg13_lv_pmos L=0.2u W=8u AS=2.12p AD=2.12p PS=13.06u
+ PD=13.06u
M$25 \$26 V\x2d \$8 \$5 sg13_lv_pmos L=0.2u W=32u AS=8.48p AD=8.48p PS=52.24u
+ PD=52.24u
M$27 \$26 V+ \$9 \$5 sg13_lv_pmos L=0.2u W=32u AS=8.48p AD=8.48p PS=52.24u
+ PD=52.24u
R$41 \$5 vdd ntap1 A=15.376p P=99.2u
R$42 \$1 gnd ptap1 A=11.376p P=75.84u
.ENDS DIFF_COMPARATOR
