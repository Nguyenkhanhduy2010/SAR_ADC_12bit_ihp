* Extracted by KLayout with SG13G2 LVS runset on : 10/02/2026 07:24

.SUBCKT C-DAC
C$1 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$2 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$3 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$4 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$5 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$6 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$7 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$8 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$9 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$10 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$11 \$7 \$4 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$12 \$7 \$4 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$13 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$14 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$15 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$16 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$17 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$18 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$19 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$20 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$21 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$22 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$23 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$24 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$25 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$26 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$27 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$28 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$29 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$30 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$31 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$32 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$33 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$34 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$35 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$36 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$37 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$38 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$39 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$40 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$41 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$42 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$43 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$44 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$45 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$46 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$47 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$48 vin|vo vref cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$49 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$50 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$51 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$52 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$53 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$54 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$55 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$56 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$57 vin|vo C4 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$58 vin|vo C4 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$59 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$60 vin|vo C1 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$61 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$62 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$63 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$64 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$65 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$66 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$67 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$68 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$69 vin|vo C4 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$70 vin|vo C3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$71 vin|vo C2 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$72 vin|vo C2 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$73 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$74 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$75 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$76 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$77 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$78 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$79 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$80 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$81 vin|vo C4 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$82 vin|vo C3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$83 vin|vo C3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$84 vin|vo C3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$85 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$86 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$87 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$88 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$89 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$90 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$91 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$92 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$93 vin|vo C4 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$94 vin|vo C4 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$95 vin|vo C4 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$96 vin|vo C4 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$97 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$98 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$99 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$100 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$101 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$102 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$103 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$104 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$105 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$106 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$107 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$108 vin|vo C5 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$109 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$110 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$111 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$112 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$113 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$114 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$115 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$116 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$117 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$118 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$119 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$120 vin|vo C6 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$121 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$122 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$123 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$124 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$125 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$126 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$127 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$128 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$129 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$130 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$131 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$132 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$133 \$5 \$3 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$134 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$135 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$136 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$137 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$138 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$139 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$140 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$141 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$142 vin|vo C_MSB cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$143 \$16 \$15 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
C$144 \$16 \$15 cap_cmim w=5.71u l=5.71u A=32.6041p P=22.84u m=1
.ENDS C-DAC
