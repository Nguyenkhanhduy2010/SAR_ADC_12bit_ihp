** sch_path: /home/designer/shared/IHP-AnalogAcademy/modules/module_3_8_bit_SAR_ADC/part_2_digital_comps/algorithm/xschem/sar_logic_tb.sch
**.subckt sar_logic_tb
V3 En GND dc 0 ac 0 PULSE(1.2 0 0 1n 1n 30u 1m)
V6 Op GND dc 0 ac 0 PULSE(1.2 0 100u 1n 1n 500u 1m)
V2 rst GND dc 0 ac 0 PULSE(0 1.2 100u 1n 1n 10u 1m)
V5 Om GND dc 0 ac 0 PULSE(0 1.2 100u 1n 1n 500u 1m)
V4 clk GND dc 0 ac 0 PULSE(0 1.2 0 10p 10p 5u 10u)
adut [ net3 net2 net4 net5 net1 ] [ net6 net7 net8 net9 net10 net11 net12 net13 net14 net15 net16 net17 net18 net19 net20 net21
+ net22 net23 net24 net25 net26 net27 ] null dut
.model dut d_cosim simulation=./sar_logic.so
A1 [ clk ] [ net3 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=0.6
A2 [ Op ] [ net2 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=0.6
A3 [ En ] [ net4 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=0.6
A4 [ Om ] [ net5 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=0.6
A5 [ rst ] [ net1 ] adc1
.model adc1 adc_bridge in_low=0.4 in_high=0.6
A6 [ net6 ] [ B5 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A7 [ net7 ] [ B4 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A8 [ net8 ] [ B3 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A9 [ net9 ] [ B2 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A10 [ net10 ] [ B1 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A11 [ net11 ] [ B0 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A12 [ net12 ] [ BN7 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A13 [ net13 ] [ BN6 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A14 [ net14 ] [ BN5 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A15 [ net15 ] [ BN4 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A16 [ net16 ] [ BN3 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A17 [ net17 ] [ BN2 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A18 [ net18 ] [ BN1 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A19 [ net19 ] [ BN0 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A20 [ net20 ] [ D7 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A21 [ net21 ] [ D6 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A22 [ net22 ] [ D5 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A23 [ net23 ] [ D4 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A24 [ net24 ] [ D3 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A25 [ net25 ] [ D2 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A26 [ net26 ] [ D1 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
A27 [ net27 ] [ D0 ] dac1
.model dac1 dac_bridge out_low=0 out_high=1.2
**** begin user architecture code


.param temp=27
.control
save all
tran 1u 200u
write sar_logic.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
