* Extracted by KLayout with SG13G2 LVS runset on : 25/02/2026 15:47

.SUBCKT bootstrap_switch gnd vdd vi vo clk
M$1 gnd clk \$3 gnd sg13_lv_nmos L=0.13u W=0.4u AS=0.136p AD=0.136p PS=1.48u
+ PD=1.48u
M$2 gnd \$3 \$4 gnd sg13_lv_nmos L=0.13u W=0.4u AS=0.136p AD=0.136p PS=1.48u
+ PD=1.48u
M$3 \$5 \$3 gnd gnd sg13_lv_nmos L=0.4u W=1.3u AS=0.442p AD=0.442p PS=3.28u
+ PD=3.28u
M$4 vi \$21 vo gnd sg13_lv_nmos L=0.13u W=2.5u AS=0.85p AD=0.85p PS=5.68u
+ PD=5.68u
M$5 \$21 vdd \$22 gnd sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$6 \$22 \$3 gnd gnd sg13_lv_nmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$7 \$5 \$7 vi gnd sg13_lv_nmos L=0.13u W=3u AS=1.02p AD=1.02p PS=6.68u PD=6.68u
M$8 gnd \$3 \$6 gnd sg13_lv_nmos L=0.13u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
M$9 \$6 vdd \$7 gnd sg13_lv_nmos L=0.13u W=3u AS=1.02p AD=1.02p PS=6.68u
+ PD=6.68u
M$10 gnd \$29 \$27 gnd sg13_lv_nmos L=0.13u W=0.4u AS=0.136p AD=0.136p PS=1.48u
+ PD=1.48u
M$11 vdd \$14 \$13 gnd sg13_lv_nmos L=0.13u W=1.3u AS=0.442p AD=0.442p PS=3.28u
+ PD=3.28u
M$12 \$14 \$13 vdd gnd sg13_lv_nmos L=0.13u W=1.3u AS=0.442p AD=0.442p PS=3.28u
+ PD=3.28u
M$13 vdd \$13 \$15 gnd sg13_lv_nmos L=0.13u W=1.3u AS=0.442p AD=0.442p PS=3.28u
+ PD=3.28u
M$14 vdd clk \$3 vdd sg13_lv_pmos L=0.13u W=0.8u AS=0.272p AD=0.272p PS=2.28u
+ PD=2.28u
M$15 vdd \$3 \$4 vdd sg13_lv_pmos L=0.13u W=0.8u AS=0.272p AD=0.272p PS=2.28u
+ PD=2.28u
M$16 \$7 \$29 vdd vdd sg13_lv_pmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$17 \$15 \$27 \$21 \$15 sg13_lv_pmos L=0.13u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$18 vdd \$29 \$27 vdd sg13_lv_pmos L=0.13u W=0.8u AS=0.272p AD=0.272p PS=2.28u
+ PD=2.28u
C$19 \$13 \$3 cap_cmim w=4.665u l=6.99u A=32.60835p P=23.31u m=1
C$20 \$14 \$4 cap_cmim w=4.665u l=6.99u A=32.60835p P=23.31u m=1
C$21 \$15 \$5 cap_cmim w=9.39u l=6.99u A=65.6361p P=32.76u m=1
.ENDS bootstrap_switch
