* Extracted by KLayout with SG13G2 LVS runset on : 14/02/2026 06:00

.SUBCKT switch_array gnd S_MSB S6 S5 S4 S3 S2 S1 D_MSB D6 D5 D4 D3 D2 D1 vref
+ \!Control|Control|vo \!Control|Control|vo$1 \!Control|Control|vo$2
+ \!Control|Control|vo$3 \!Control|Control|vo$4 \!Control|Control|vo$5 vdd
+ \!Control|Control|vo$6
M$1 vref \!Control|Control|vo$1 S6 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p
+ AD=0.34p PS=2.68u PD=2.68u
M$2 gnd D6 S6 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$3 vref \!Control|Control|vo S_MSB gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p
+ AD=0.34p PS=2.68u PD=2.68u
M$4 gnd D_MSB S_MSB gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u
+ PD=2.68u
M$5 vref \!Control|Control|vo$5 S1 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p
+ AD=0.34p PS=2.68u PD=2.68u
M$6 gnd D1 S1 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$7 vref \!Control|Control|vo$2 S5 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p
+ AD=0.34p PS=2.68u PD=2.68u
M$8 vref \!Control|Control|vo$3 S4 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p
+ AD=0.34p PS=2.68u PD=2.68u
M$9 vref \!Control|Control|vo$4 S3 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p
+ AD=0.34p PS=2.68u PD=2.68u
M$10 gnd D5 S5 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$11 gnd D4 S4 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$12 gnd D3 S3 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$13 vref \!Control|Control|vo$6 S2 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p
+ AD=0.34p PS=2.68u PD=2.68u
M$14 gnd D2 S2 gnd sg13_lv_nmos L=0.13u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$15 gnd D6 \!Control|Control|vo$1 gnd sg13_lv_nmos L=0.13u W=0.4u AS=0.136p
+ AD=0.136p PS=1.48u PD=1.48u
M$16 gnd D_MSB \!Control|Control|vo gnd sg13_lv_nmos L=0.13u W=0.4u AS=0.136p
+ AD=0.136p PS=1.48u PD=1.48u
M$17 gnd D1 \!Control|Control|vo$5 gnd sg13_lv_nmos L=0.13u W=0.4u AS=0.136p
+ AD=0.136p PS=1.48u PD=1.48u
M$18 gnd D5 \!Control|Control|vo$2 gnd sg13_lv_nmos L=0.13u W=0.4u AS=0.136p
+ AD=0.136p PS=1.48u PD=1.48u
M$19 gnd D4 \!Control|Control|vo$3 gnd sg13_lv_nmos L=0.13u W=0.4u AS=0.136p
+ AD=0.136p PS=1.48u PD=1.48u
M$20 gnd D3 \!Control|Control|vo$4 gnd sg13_lv_nmos L=0.13u W=0.4u AS=0.136p
+ AD=0.136p PS=1.48u PD=1.48u
M$21 gnd D2 \!Control|Control|vo$6 gnd sg13_lv_nmos L=0.13u W=0.4u AS=0.136p
+ AD=0.136p PS=1.48u PD=1.48u
M$22 vdd D6 \!Control|Control|vo$1 vdd sg13_lv_pmos L=0.13u W=0.8u AS=0.272p
+ AD=0.272p PS=2.28u PD=2.28u
M$23 vdd D_MSB \!Control|Control|vo vdd sg13_lv_pmos L=0.13u W=0.8u AS=0.272p
+ AD=0.272p PS=2.28u PD=2.28u
M$24 vdd D1 \!Control|Control|vo$5 vdd sg13_lv_pmos L=0.13u W=0.8u AS=0.272p
+ AD=0.272p PS=2.28u PD=2.28u
M$25 vdd D5 \!Control|Control|vo$2 vdd sg13_lv_pmos L=0.13u W=0.8u AS=0.272p
+ AD=0.272p PS=2.28u PD=2.28u
M$26 vdd D4 \!Control|Control|vo$3 vdd sg13_lv_pmos L=0.13u W=0.8u AS=0.272p
+ AD=0.272p PS=2.28u PD=2.28u
M$27 vdd D3 \!Control|Control|vo$4 vdd sg13_lv_pmos L=0.13u W=0.8u AS=0.272p
+ AD=0.272p PS=2.28u PD=2.28u
M$28 vdd D2 \!Control|Control|vo$6 vdd sg13_lv_pmos L=0.13u W=0.8u AS=0.272p
+ AD=0.272p PS=2.28u PD=2.28u
M$29 vref D6 S6 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
M$30 gnd \!Control|Control|vo$1 S6 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p
+ AD=0.68p PS=4.68u PD=4.68u
M$31 vref D_MSB S_MSB vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
M$32 gnd \!Control|Control|vo S_MSB vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p
+ AD=0.68p PS=4.68u PD=4.68u
M$33 vref D1 S1 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
M$34 gnd \!Control|Control|vo$5 S1 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p
+ AD=0.68p PS=4.68u PD=4.68u
M$35 vref D5 S5 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
M$36 vref D4 S4 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
M$37 vref D3 S3 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
M$38 gnd \!Control|Control|vo$2 S5 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p
+ AD=0.68p PS=4.68u PD=4.68u
M$39 gnd \!Control|Control|vo$3 S4 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p
+ AD=0.68p PS=4.68u PD=4.68u
M$40 gnd \!Control|Control|vo$4 S3 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p
+ AD=0.68p PS=4.68u PD=4.68u
M$41 vref D2 S2 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
M$42 gnd \!Control|Control|vo$6 S2 vdd sg13_lv_pmos L=0.13u W=2u AS=0.68p
+ AD=0.68p PS=4.68u PD=4.68u
.ENDS switch_array
